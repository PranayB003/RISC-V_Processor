`define WORD_WIDTH     32
`define REG_ADDR_WIDTH 5
`define IMEM_DEPTH     1024
`define DMEM_DEPTH     1024
