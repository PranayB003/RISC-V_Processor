`define WORDSZ    32
`define NREGS     32
`define REGADDRSZ 5
`define IMEMSZ    1024
`define DMEMSZ    1024
